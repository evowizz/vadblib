// Copyright 2023 Dylan Roussel
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
module vadblib

[params]
pub struct StartRestartParams {
	port u16 = 5037
}

// start runs the command `adb -P {port} start-server` where `{port}`
// is provided with the optional parameter `params.port`.
pub fn (adb AndroidDebugBridge) start(params StartRestartParams) ! {
	adb.run(command: '-P ${params.port} start-server')!
}

// kill runs the command `adb kill-server`.
pub fn (adb AndroidDebugBridge) kill() ! {
	adb.run(command: 'kill-server')!
}

// restart runs the commands `adb kill-server` followed by
// `adb -P {port} start-server` where `{port}` is provided with
// the optional parameter `params.port`.
pub fn (adb AndroidDebugBridge) restart(params StartRestartParams) ! {
	adb.kill()!
	adb.start(params)!
}
